
// ====================================================================================================
// ====================================================================================================

shift( dir ,
       val ,
       in  ,
       out );

endmodule: shift

// ====================================================================================================
// ====================================================================================================

module sctrl(
    opcode ,
    sdiff  ,
    s1     ,
    s2     ,
    inv1   ,
    inv2
);

// --------------------------------------------------
parameter S = 1 ;
parameter E = 8 ;
parameter M = 23;

// --------------------------------------------------
input   opcode  ;
input   sdiff   ;
input   s1      ;
input   s2      ;

output  inv1    ;
output  inv2    ;

// --------------------------------------------------

endmodule: sctrl

// ====================================================================================================
// ====================================================================================================

module adder( a ,
              b ,
              c );

// --------------------------------------------------
parameter S = 1 ;
parameter E = 8 ;
parameter M = 23;

// --------------------------------------------------
input    [M-1:0] a;
input    [M-1:0] b;
output   [M-1:0] c;

// --------------------------------------------------

endmodule: adder

// ====================================================================================================
// ====================================================================================================

module complement(
    in,
    out,
    enable
);

// --------------------------------------------------
parameter S = 1 ;
parameter E = 8 ;
parameter M = 23;

// --------------------------------------------------
input               enable ;
input   [M-1:0]     in     ;
output  [M-1:0]     out    ;

// --------------------------------------------------
wire              enable ;
wire  [M-1:0]     in     ;
wire  [M-1:0]     out    ;

// --------------------------------------------------
assign out[M-1:0] = (enable) ? (~in[M-1:0] + 1'b1) : in[M-1:0];

endmodule:complement

// ====================================================================================================
// Opcode : Add=0 ; Sub=1 ;
// ====================================================================================================

module fpu(
    operand1 ,
    operand2 ,
    opcode   ,
    result   
    );

// --------------------------------------------------
parameter S = 1 ;
parameter E = 8 ;
parameter M = 23;

// --------------------------------------------------
// InOut
input               opcode ;
input  [S+E+M-1:0]  op1    ;
input  [S+E+M-1:0]  op2    ;
output [S+E+M-1:0]  result ;

wire              opcode ;
wire [S+E+M-1:0]  op1    ;
wire [S+E+M-1:0]  op2    ;
wire [S+E+M-1:0]  result ;

// --------------------------------------------------
// Wiring



// --------------------------------------------------
// Instances

// COMP

// SCTRL
sctrl #( .S(S), .E(E), .M(M)) fpu_sctrl (
    // In
    .opcode ( opcode ) ,
    .sdiff  ( sdiff  ) ,
    .s1     ( s1     ) ,
    .s2     ( s2     ) ,
    // Out
    .inv1   ( inv1   ) ,
    .inv2   ( inv2   ) ,
    );

// 1st Level
wire [M-1:0]    m1;
wire [M-1:0]    m2;

wire [M-1:0]    m1_muxed;
wire [M-1:0]    m2_muxed;

assign m1_muxed = (sdiff) ? m1 : m2;
assign m2_muxed = (sdiff) ? m2 : m1;

// RShift
rshift #( .S(S), .E(E), .M(M)) fpu_rshift (
    .dir ( 0          ) , // right=0 left=1
    .val ( rshift_val ) ,
    .in  ( m2_muxed   ) ,
    .out ( rshift_out )
    );

// Complements
complement #( .S(S), .E(E), .M(M)) m1_complement (
    .enable ( inv1              ) ,
    .in     ( m1_muxed          ) ,
    .out    ( m1_complement_out )
);

complement #( .S(S), .E(E), .M(M)) m2_complement (
    .enable ( inv2              ) ,
    .in     ( rshift_out        ) ,
    .out    ( m2_complement_out )
);

endmodule: fpu



